library verilog;
use verilog.vl_types.all;
entity micro_tb_v is
end micro_tb_v;
