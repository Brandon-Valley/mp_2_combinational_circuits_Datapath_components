library verilog;
use verilog.vl_types.all;
entity deMUX_1_8_tb_v is
end deMUX_1_8_tb_v;
