library verilog;
use verilog.vl_types.all;
entity priority_enc_4_2_tb_v is
end priority_enc_4_2_tb_v;
