library verilog;
use verilog.vl_types.all;
entity \OR4_v__equation\ is
    port(
        i_a             : in     vl_logic;
        i_b             : in     vl_logic;
        i_c             : in     vl_logic;
        i_d             : in     vl_logic;
        o_f             : out    vl_logic
    );
end \OR4_v__equation\;
