library verilog;
use verilog.vl_types.all;
entity SN74145_tb_v is
end SN74145_tb_v;
