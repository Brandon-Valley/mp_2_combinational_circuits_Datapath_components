library verilog;
use verilog.vl_types.all;
entity MUX_4_1_8_bit_tb_v is
end MUX_4_1_8_bit_tb_v;
