// -- python C:\Users\Brandon\Documents\Personal_Projects\my_utils\modelsim_utils\auto_run.py -d run_cmd__XOR4_v.do

////////////////////////////////
// Equation Model
////////////////////////////////
module XOR4_v__equation
  (input i_a, i_b, i_c, i_d,
   output o_f);
   
  assign o_f = (i_a ^ i_b) ^ (i_c ^ i_d);
  
endmodule


////////////////////////////////
// Behavior Model
////////////////////////////////
module XOR4_v__behavior
  (input i_a, i_b, i_c, i_d,
   output o_f);
   
  assign o_f = (~ i_a & ~ i_b & ~ i_c &   i_d) | 
               (~ i_a & ~ i_b &   i_c & ~ i_d) |
               (~ i_a &   i_b & ~ i_c & ~ i_d) |
               (  i_a & ~ i_b & ~ i_c & ~ i_d) |
               (  i_a &   i_b &   i_c & ~ i_d) |
               (  i_a &   i_b & ~ i_c &   i_d) |
               (  i_a & ~ i_b &   i_c &   i_d) |
               (~ i_a &   i_b &   i_c &   i_d) ? 1 : 0;
  
endmodule



////////////////////////////////
// Component Model - Self
////////////////////////////////
module XOR4_v__cmpnt_self
  (input i_a, i_b, i_c, i_d,
  output o_f);
   
  wire fi1, fi2; // internal outputs
   
  XOR2_v xor1 (i_a, i_b, fi1);
  XOR2_v xor2 (i_c, i_d, fi2);
  XOR2_v xor3 (fi1, fi2, o_f);

    
endmodule


// ////////////////////////////////
// // Component Model - Primative
// ////////////////////////////////
// module XOR4_v__cmpnt_prim
  // (input i_a, i_b, i_c, i_d,
  // output o_f);
   
  // wire fi1, fi2, fi3; // internal outputs
   
  // AND2_v and1 (i_a, i_b, fi1);
  // AND2_v and2 (i_c, i_d, fi2);
  // AND2_v and3 (fi1, fi2, fi3);
  // NOT1_v not1 (fi3, o_f);

    
// endmodule





