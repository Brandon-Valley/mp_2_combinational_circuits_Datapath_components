library verilog;
use verilog.vl_types.all;
entity priority_enc_8_3_tb_v is
end priority_enc_8_3_tb_v;
