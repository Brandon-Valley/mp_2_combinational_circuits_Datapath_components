library verilog;
use verilog.vl_types.all;
entity NAND4_tb_v is
end NAND4_tb_v;
