library verilog;
use verilog.vl_types.all;
entity XOR4_tb_v is
end XOR4_tb_v;
