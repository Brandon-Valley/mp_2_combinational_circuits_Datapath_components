library verilog;
use verilog.vl_types.all;
entity MUX_8_1_tb_v is
end MUX_8_1_tb_v;
