library verilog;
use verilog.vl_types.all;
entity OR4_tb_v_TEST is
end OR4_tb_v_TEST;
