library verilog;
use verilog.vl_types.all;
entity MUX_4_1_2_bit_tb_v is
end MUX_4_1_2_bit_tb_v;
