library verilog;
use verilog.vl_types.all;
entity NOT1_v is
    port(
        i_a             : in     vl_logic;
        o_f             : out    vl_logic
    );
end NOT1_v;
